module four_bit_RCA_RCS(A, B, Cin, S, Cout);
input [3:0] A, B;
input Cin;
output [3:0] S;
output Cout;
wire c1, c2, c3;
one_bit_full_adder FA0(A[0], B[0], Cin, S[0], c1);
one_bit_full_adder FA1(A[1], B[1], c1, S[1], c2);
one_bit_full_adder FA2(A[2], B[2], c2, S[2], c3);
one_bit_full_adder FA3(A[3], B[3], c3, S[3], Cout);
endmodule

module one_bit_full_adder(A, B, Cin, S, Cout);
input A, B, Cin;
output S, Cout;
wire and_0_out, and_1_out, and_2_out, xor_0_out;
xor (xor_0_out, A, B);
xor (S, xor_0_out, Cin);
and (and_0_out, A, B);
and (and_1_out, B, Cin);
and (and_2_out, A, Cin);
or (Cout, and_0_out, and_1_out, and_2_out);
endmodule

module CLA(A, B, Cin, S, Cout);
input [31:0] A, B;
input Cin;
output [31:0] S;
output Cout;
wire [7:0] P, G;
wire [8:0] C;
assign C[0] = Cin;
assign Cout = C[8];
wire [7:0] block_cout;
four_bit_RCA_RCS RCA0(A[3:0], B[3:0], C[0], S[3:0], block_cout[0]);
four_bit_RCA_RCS RCA1(A[7:4], B[7:4], C[1], S[7:4], block_cout[1]);
four_bit_RCA_RCS RCA2(A[11:8], B[11:8], C[2], S[11:8], block_cout[2]);
four_bit_RCA_RCS RCA3(A[15:12], B[15:12], C[3], S[15:12], block_cout[3]);
four_bit_RCA_RCS RCA4(A[19:16], B[19:16], C[4], S[19:16], block_cout[4]);
four_bit_RCA_RCS RCA5(A[23:20], B[23:20], C[5], S[23:20], block_cout[5]);
four_bit_RCA_RCS RCA6(A[27:24], B[27:24], C[6], S[27:24], block_cout[6]);
four_bit_RCA_RCS RCA7(A[31:28], B[31:28], C[7], S[31:28], block_cout[7]);
wire p0, p1, p2, p3, g0, g1, g2, g3;
assign p0 = A[0] | B[0];
assign p1 = A[1] | B[1];
assign p2 = A[2] | B[2];
assign p3 = A[3] | B[3];
assign g0 = A[0] & B[0];
assign g1 = A[1] & B[1];
assign g2 = A[2] & B[2];
assign g3 = A[3] & B[3];
assign P[0] = p0 & p1 & p2 & p3;
assign G[0] = g3 | (p3 & g2) | (p3 & p2 & g1) | (p3 & p2 & p1 & g0);
wire p4, p5, p6, p7, g4, g5, g6, g7;
assign p4 = A[4] | B[4];
assign p5 = A[5] | B[5];
assign p6 = A[6] | B[6];
assign p7 = A[7] | B[7];
assign g4 = A[4] & B[4];
assign g5 = A[5] & B[5];
assign g6 = A[6] & B[6];
assign g7 = A[7] & B[7];
assign P[1] = p4 & p5 & p6 & p7;
assign G[1] = g7 | (p7 & g6) | (p7 & p6 & g5) | (p7 & p6 & p5 & g4);
wire p8, p9, p10, p11, g8, g9, g10, g11;
assign p8 = A[8] | B[8];
assign p9 = A[9] | B[9];
assign p10 = A[10] | B[10];
assign p11 = A[11] | B[11];
assign g8 = A[8] & B[8];
assign g9 = A[9] & B[9];
assign g10 = A[10] & B[10];
assign g11 = A[11] & B[11];
assign P[2] = p8 & p9 & p10 & p11;
assign G[2] = g11 | (p11 & g10) | (p11 & p10 & g9) | (p11 & p10 & p9 & g8);
wire p12, p13, p14, p15, g12, g13, g14, g15;
assign p12 = A[12] | B[12];
assign p13 = A[13] | B[13];
assign p14 = A[14] | B[14];
assign p15 = A[15] | B[15];
assign g12 = A[12] & B[12];
assign g13 = A[13] & B[13];
assign g14 = A[14] & B[14];
assign g15 = A[15] & B[15];
assign P[3] = p12 & p13 & p14 & p15;
assign G[3] = g15 | (p15 & g14) | (p15 & p14 & g13) | (p15 & p14 & p13 & g12);
wire p16, p17, p18, p19, g16, g17, g18, g19;
assign p16 = A[16] | B[16];
assign p17 = A[17] | B[17];
assign p18 = A[18] | B[18];
assign p19 = A[19] | B[19];
assign g16 = A[16] & B[16];
assign g17 = A[17] & B[17];
assign g18 = A[18] & B[18];
assign g19 = A[19] & B[19];
assign P[4] = p16 & p17 & p18 & p19;
assign G[4] = g19 | (p19 & g18) | (p19 & p18 & g17) | (p19 & p18 & p17 & g16);
wire p20, p21, p22, p23, g20, g21, g22, g23;
assign p20 = A[20] | B[20];
assign p21 = A[21] | B[21];
assign p22 = A[22] | B[22];
assign p23 = A[23] | B[23];
assign g20 = A[20] & B[20];
assign g21 = A[21] & B[21];
assign g22 = A[22] & B[22];
assign g23 = A[23] & B[23];
assign P[5] = p20 & p21 & p22 & p23;
assign G[5] = g23 | (p23 & g22) | (p23 & p22 & g21) | (p23 & p22 & p21 & g20);
wire p24, p25, p26, p27, g24, g25, g26, g27;
assign p24 = A[24] | B[24];
assign p25 = A[25] | B[25];
assign p26 = A[26] | B[26];
assign p27 = A[27] | B[27];
assign g24 = A[24] & B[24];
assign g25 = A[25] & B[25];
assign g26 = A[26] & B[26];
assign g27 = A[27] & B[27];
assign P[6] = p24 & p25 & p26 & p27;
assign G[6] = g27 | (p27 & g26) | (p27 & p26 & g25) | (p27 & p26 & p25 & g24);
wire p28, p29, p30, p31, g28, g29, g30, g31;
assign p28 = A[28] | B[28];
assign p29 = A[29] | B[29];
assign p30 = A[30] | B[30];
assign p31 = A[31] | B[31];
assign g28 = A[28] & B[28];
assign g29 = A[29] & B[29];
assign g30 = A[30] & B[30];
assign g31 = A[31] & B[31];
assign P[7] = p28 & p29 & p30 & p31;
assign G[7] = g31 | (p31 & g30) | (p31 & p30 & g29) | (p31 & p30 & p29 & g28);
assign C[1] = G[0] | (P[0] & C[0]);
assign C[2] = G[1] | (P[1] & C[1]);
assign C[3] = G[2] | (P[2] & C[2]);
assign C[4] = G[3] | (P[3] & C[3]);
assign C[5] = G[4] | (P[4] & C[4]);
assign C[6] = G[5] | (P[5] & C[5]);
assign C[7] = G[6] | (P[6] & C[6]);
assign C[8] = G[7] | (P[7] & C[7]);
endmodule
